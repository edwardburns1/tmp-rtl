// Code your testbench here


//`include "top_testbench.sv"
//`include "PC_testbench.sv"
//`include "reg_file_testbench.sv"

//`include "ALU_testbench.sv"
`include "top_testbench.sv"