// Code your design here
`include "PC.sv"
`include "reg_file.sv"
`include "ALU.sv"