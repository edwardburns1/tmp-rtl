// Code your design here
`include "PC.sv"
`include "reg_file.sv"
`include "ALU.sv"
`include "fetch.sv"
`include "decode_execute.sv"
`include "write_back.sv"
`include "top_level.sv"