module write_back(
    input wire clk,           
    input wire reset,            
    input wire [31:0] result,  
    input write_enable,
    input wire  [31:0] write address
);

  
  //if write enable then write back to the register? 


endmodule