module write_back(
    input wire clk,           
    input wire reset,      
    inout wire [31:0] memory [0:1023], // Memory input
    input wire [31:0] result,  
    input reg_write_enable
  //input wire  [31:0] store_memory_address
  //
);

  
  //if write enable then write back to the register? 
  /*
   if (reg_write_enable)
   	
  */


endmodule